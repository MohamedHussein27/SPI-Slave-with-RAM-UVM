package spi_slave_driver_pkg;
    import spi_slave_shared_pkg::*;
    import spi_slave_config_obj_pkg::*;
    import spi_slave_seq_item_pkg::*;
    import uvm_pkg::*;
    `include "uvm_macros.svh"    
    class spi_slave_driver extends uvm_driver #(spi_slave_seq_item);
        `uvm_component_utils(spi_slave_driver)

        virtual spi_slave_if spi_slave_vif; // virtual interface
        spi_slave_seq_item stim_seq_item; // sequence item

        function new(string name = "spi_slave_driver", uvm_component parent = null);
            super.new(name, parent);
        endfunction

        task run_phase(uvm_phase phase);
            super.run_phase(phase);
            forever begin
                stim_seq_item = spi_slave_seq_item::type_id::create("stim_seq_item");
                seq_item_port.get_next_item(stim_seq_item);
                spi_slave_vif.rst_n = stim_seq_item.rst_n;
                spi_slave_vif.MOSI = stim_seq_item.MOSI;
                sampling_MOSI = stim_seq_item.MOSI;
                spi_slave_vif.tx_valid = stim_seq_item.tx_valid;
                spi_slave_vif.ss_n = stim_seq_item.ss_n;
                spi_slave_vif.tx_data = stim_seq_item.tx_data;
                #20;
                seq_item_port.item_done();
                `uvm_info("run_phase", stim_seq_item.convert2string_stimulus(), UVM_HIGH)
            end
        endtask
    endclass
endpackage
            
