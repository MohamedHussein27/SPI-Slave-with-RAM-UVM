package spi_slave_shared_pkg;
    typedef enum {IDLE, CHK_CMD, WRITE, READ_ADD, READ_DATA} cs_e;
    cs_e cs; // i defined cs here so it can be accessed by both scoreboard and testbench
    cs_e ns; // next state logic
    // internal signals
    int counter = 0; // counter used in reference model in READ_DATA state to verify MISO_ref Correctly
    bit state_finished; // when high, that means the current state is finished 
    bit tx_flag = 0; // flag to make tx_valid high while READ_DATA state
    bit delay; // just a falg to add 1 clock delay to synchronize between dut and reference model
    int i; // counter used in reaad_add constriant
    bit write_constraint; // flag to lock and open write constraints on MOSI
    bit read_add_constraint; // flag to lock and open read address constraints on MOSI
    bit read_data_constraint; // flag to lock and open read data constraints on MOSI
    // counters
    int correct_count_out = 0;
    int error_count_out = 0;
endpackage
