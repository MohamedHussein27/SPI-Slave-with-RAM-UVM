package ram_shared_pkg;
    int error_count_out = 0; 
    int correct_count_out = 0;
endpackage